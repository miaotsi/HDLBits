module top_module( 
    input in, 
    output out 
);
	
    //assign out = ~in; //按照位非
    assign out = !in;　// 逻辑非

endmodule
